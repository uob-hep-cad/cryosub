.title KiCad schematic
.include "/Users/phdgc/Downloads/MMBFJ201.lib"
R4 Net-_Q1-Pad2_ 0 1.5k
V1 VDD 0 dc 10
JQ1 VDD Net-_Q1-Pad2_ 0 MMBFJ201
.end
