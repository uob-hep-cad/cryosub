.title KiCad schematic
.include "../FDD306P.lib"
XQ1 /vload /vcont /vdd FDD306P
V1 /vdd 0 dc 5
V2 /vcont 0 pulse(0 5 0 10 10 20 40)
R1 /vload 0 5
.end
