.title KiCad schematic
.include "./IFX-Power_OptiMOS_N-channel_small_signal_MOSFET_240V_250V_400V_600V_Spice-web.lib"
R7 Net-_R6-Pad2_ 0 30k
V2 /vg2 Net-_R6-Pad2_ dc 0 ac 1 sin(0 500m 1k)
R6 VDD Net-_R6-Pad2_ 20k
XQ2 /vd2 /vg2 /vs BSS127_L0
V1 VDD 0 dc 5
XQ1 /vd1 /vg1 /vs BSS127_L0
R5 VDD /vd2 4.7k
R9 /vg1 /vd2 200k
R3 VDD /vd1 4.7k
R8 /vd1 /vg2 200k
R1 VDD /vg1 20k
R4 /vs 0 1K
R2 /vg1 0 30k
.TEMP 27 
.CONTROL ABSTOL=1nA CHGTOL=1pC ITL1=150 ITL2=150 ITL4=500 RELTOL=0.011 
.ENDC 
.IC V(/vd1 )=4.5  V(/vd2)=2.0 
.end
