.title KiCad schematic
.include "./FDD306P.lib"
.include "./IFX-Power_OptiMOS_N-channel_small_signal_MOSFET_240V_250V_400V_600V_Spice-web.lib"
.include "./sim_ntc_10k_1.lib"
.include "RB751V40T1G.lib"
R7 5V0 /vg2 6.8k
V2 /vtemp 0 dc 270 ac 1 pulse(1 350 0 10 10 10 100)
XQ2 /vd2 /vg2 /vs BSS127_L0
V1 5V0 0 dc 5
XQ1 /vd1 /vg1 /vs BSS127_L0
R5 5V0 /vd2 4.7k
R9 /vg1 /vd2 20k
R3 5V0 /vd1 4.7k
R8 /vd1 /vg2 20k
R1 5V0 /vg1 6.8k
R4 /vs 0 1K
R2 /vg1 0 10k
XTH1 /vg2 0 /vtemp 0 NTC_10K_1
XQ3 /vload /vg3 5V0 FDD306P
R6 /vload 0 5
C2 /vload 0 1u
C1 /vload /vg3 30n
R10 /vg3 Net-_D1-Pad1_ 1k
D1 /vd2 Net-_D1-Pad1_ rb751v40t1g
R11 /vg3 0 100k
R12 /vg3 Net-_D2-Pad1_ 1k
D2 0 Net-_D2-Pad1_ rb751v40t1g
.TEMP 27 
.CONTROL 
OPTIONS ABSTOL=1nA CHGTOL=1pC ITL1=150 ITL2=150 ITL4=500 RELTOL=0.011
tran 5m 30
set filetype=ascii 
set wr_vecnames 
set wr_singlescale 
wrdata tmp.txt V( "/vd1" ) V("/vd2") V("/vtemp") V("/vload") 
.ENDC 
.end
